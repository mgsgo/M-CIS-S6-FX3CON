# This file was generated with hex2rom written by Daniel Wallner

INST *brom231300 INIT_00 = 1D01B0A010D1B1A00D31C803F1E8B0A010CDCF1F111A1B1C1D1E1F202122230A;
INST *brom231300 INIT_01 = E008D0C01908F7E6DFCF1F0FFFEF088CFE5F08899A98088CFE5DDA7559E1B1A1;
INST *brom231300 INIT_02 = 06DFCEF9FDECDFCEE8DFCF1F0FFFEF08EFFF0F1FCFDFACDFCE21E0901F0E81F1;
INST *brom231300 INIT_03 = 82818F08EFFF0F1FCFDF618888FDEC09F1E0908D298A80FFEE2109F1E0900F10;
INST *brom231300 INIT_04 = 4120534DFFF8F29695A980F7961189FB951188A1C59086A970659080898A8A88;
INST *brom231300 INIT_05 = 0000000000000000000000000000000000000000007374656F20667333335339;
INST *brom231301 INIT_00 = 92C0E0E8E0F70738929695C0E0E3E0E6E0BFEDBE24C0C0C0C0C0C0C0C0C0C0C0;
INST *brom231301 INIT_01 = 2FC0E0E02F2F2E2E93939393929295B1CF9B95B9B9E195B9CF9BCFC0D0F70738;
INST *brom231301 INIT_02 = E22D2D2E2E2E2D2D2E93939393929295909091919191F3051596DFE02F2F912F;
INST *brom231301 INIT_03 = BBBBEF95909091919191F723812E2E952F2FE0E0F430812D2D96952F2FE0C0E0;
INST *brom231301 INIT_04 = 54004747CF94CF9898F733CF9AF433CF9AF433DFDFE0E6DFE0E0E0E6B9E1B9E1;
INST *brom231301 INIT_05 = 0000000000000000000000000000000000000000007465207263746F20313230;
