-- $Id: mem1.vhd,v 1.2 2008/05/27 18:57:39 jrothwei Exp jrothwei $
-- Joseph Rothweiler, Sensicomm LLC, Started 21May2008.
--
-- Copyright 2008 Sensicomm LLC
--
-- This program is free software: you can redistribute it and/or modify
-- it under the terms of the GNU General Public License as published by
-- the Free Software Foundation, either version 3 of the License, or
-- (at your option) any later version.
--
-- This program is distributed in the hope that it will be useful,
-- but WITHOUT ANY WARRANTY; without even the implied warranty of
-- MERCHANTABILITY or FITNESS FOR A PARTICULAR PURPOSE.  See the
-- GNU General Public License for more details.
--
-- You should have received a copy of the GNU General Public License
-- along with this program.  If not, see <http://www.gnu.org/licenses/>.

-- Testing the AX8 core from opencores.org, which implements
-- most of the Atmel AVR instruction set. This top-level file
-- is loosely based on the A90S2313 file from the AX8 package,
-- but it is no longer attempting to copy a specific Atmel chip.
-- A Xilinx RAM block is now used for program memory, so it can
-- be updated.

-- Creating a 1kx16 RAM block for use by the AX8 core.
----------------------------------------------------------------------------------
library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

library UNISIM;
use UNISIM.VComponents.all;

entity mem_1kx16 is
    Port ( Clk : in  STD_LOGIC;
           A : in  STD_LOGIC_VECTOR(9 downto 0);   -- Address
           D : out  STD_LOGIC_VECTOR(15 downto 0)  -- Data_out
    );
end mem_1kx16;

architecture Behavioral of mem_1kx16 is
   -- These are dummy signals, for memory ports that aren't currently used.
   signal DOA : STD_LOGIC_VECTOR(16-1 downto 0);
   signal DOB : STD_LOGIC_VECTOR(7 downto 0);
   signal DOPA : STD_LOGIC_VECTOR(1 downto 0);
   signal DOPB : STD_LOGIC_VECTOR(0 downto 0); -- Does this work???
   signal ADDRB : STD_LOGIC_VECTOR(10 downto 0) := "000" & X"00"; 
   signal CLKB : STD_LOGIC := '1';
   signal DIA : STD_LOGIC_VECTOR(15 downto 0) := X"FFFF";
   signal DIB : STD_LOGIC_VECTOR(7 downto 0) := X"FF";
   signal DIPA : STD_LOGIC_VECTOR(1 downto 0) := "11";
   signal DIPB : STD_LOGIC_VECTOR(0 downto 0) := "1" ; -- Does this work???
   signal ENA : STD_LOGIC := '0';  -- Enable port A
   signal ENB : STD_LOGIC := '0';  -- Disable port B for now.
   signal SSRA : STD_LOGIC := '0'; -- Don't use the output resets.
   signal SSRB : STD_LOGIC := '0'; -- Don't use the output resets.
   signal WEA : STD_LOGIC_VECTOR(1 downto 0) := "00"; -- No writes at all for now.
   signal WEB : STD_LOGIC := '0'; -- No writes at all for now.

begin

	ADDRB		<= '0' & A;

   -- RAMB16BWE_S18_S9: 1k/2k x 16/8 + 2/1 Parity bits Dual-Port byte-wide write RAM
   --                   Spartan-3A 
   -- Xilinx HDL Language Template, version 10.1.1

   RAMB16BWE_S18_S9_inst_LSB : RAMB16BWE_S18_S9
   generic map (
      INIT_A => X"00000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      SRVAL_A => X"00000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      -- The following INIT_xx declarations specify the intiial contents of the RAM
      -- Port A Address 0 to 255, Port B address 0 to 127
      --INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Program pgm_blink.asm, manually entered
      --           .   .   .   .   .   .   .   .   .   .   .   .   .   .   .   .
      INIT_00 => X"1D01B0A010D1B1A00D31C803F1E8B0A010CDCF1F111A1B1C1D1E1F202122230A",
      INIT_01 => X"E008D0C01908F7E6DFCF1F0FFFEF088CFE5F08899A98088CFE5DDA7559E1B1A1",
      INIT_02 => X"06DFCEF9FDECDFCEE8DFCF1F0FFFEF08EFFF0F1FCFDFACDFCE21E0901F0E81F1",
      INIT_03 => X"82818F08EFFF0F1FCFDF618888FDEC09F1E0908D298A80FFEE2109F1E0900F10",
      INIT_04 => X"4120534DFFF8F29695A980F7961189FB951188A1C59086A970659080898A8A88",
      INIT_05 => X"0000000000000000000000000000000000000000007374656F20667333335339",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 256 to 511, Port B Address 128 to 255
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 512 to 767, Port B Address 256 to 383
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 768 to 1023, Port B Address 384 to 511
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Port A Address 0 to 255, Port B Address 0 to 127
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 256 to 511, Port B Address 128 to 255
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 512 to 767, Port B Address 256 to 383
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 768 to 1023, Port B Address 384 to 511
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => open,--DOA,    --  DOA,      -- Port A 16-bit Data Output
      DOB => D(8-1 downto 0),--D(16-1 downto 8),--DOB,      -- Port B 8-bit Data Output
      DOPA => open,--DOPA,    -- Port A 2-bit Parity Output
      DOPB => open,--DOPB,    -- Port B 1-bit Parity Output
      ADDRA => "0000000000",--A,  --  ADDRA,  -- Port A 10-bit Address Input
      ADDRB => ADDRB,  -- Port B 11-bit Address Input
      CLKA => '0',--Clk, --  CLKA,    -- Port A 1-bit Clock
      CLKB => Clk,--CLKB,    -- Port B 1-bit Clock
      DIA => DIA,      -- Port A 16-bit Data Input
      DIB => DIB,      -- Port B 8-bit Data Input
      DIPA => DIPA,    -- Port A 2-bit parity Input
      DIPB => DIPB,    -- Port B 1-bit parity Input
      ENA => ENA,      -- Port A 1-bit RAM Enable Input
      ENB => '1',--ENB,      -- Port B 1-bit RAM Enable Input
      SSRA => SSRA,    -- Port A 1-bit Synchronous Set/Reset Input
      SSRB => SSRB,    -- Port B 1-bit Synchronous Set/Reset Input
      WEA => WEA,      -- Port A 2-bit Write Enable Input
      WEB => WEB       -- Port B 1-bit Write Enable Input
   );

   RAMB16BWE_S18_S9_inst_MSB : RAMB16BWE_S18_S9
   generic map (
      INIT_A => X"00000", --  Value of output RAM registers on Port A at startup
      INIT_B => X"000", --  Value of output RAM registers on Port B at startup
      SIM_COLLISION_CHECK => "ALL", -- "NONE", "WARNING", "GENERATE_X_ONLY", "ALL" 
      SRVAL_A => X"00000", --  Port A ouput value upon SSR assertion
      SRVAL_B => X"000", --  Port B ouput value upon SSR assertion
      WRITE_MODE_A => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      WRITE_MODE_B => "READ_FIRST", --  WRITE_FIRST, READ_FIRST or NO_CHANGE
      -- The following INIT_xx declarations specify the intiial contents of the RAM
      -- Port A Address 0 to 255, Port B address 0 to 127
      --INIT_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Program pgm_blink.asm, manually entered
      --           .   .   .   .   .   .   .   .   .   .   .   .   .   .   .   .
      INIT_00 => X"92C0E0E8E0F70738929695C0E0E3E0E6E0BFEDBE24C0C0C0C0C0C0C0C0C0C0C0",
      INIT_01 => X"2FC0E0E02F2F2E2E93939393929295B1CF9B95B9B9E195B9CF9BCFC0D0F70738",
      INIT_02 => X"E22D2D2E2E2E2D2D2E93939393929295909091919191F3051596DFE02F2F912F",
      INIT_03 => X"BBBBEF95909091919191F723812E2E952F2FE0E0F430812D2D96952F2FE0C0E0",
      INIT_04 => X"54004747CF94CF9898F733CF9AF433CF9AF433DFDFE0E6DFE0E0E0E6B9E1B9E1",
      INIT_05 => X"0000000000000000000000000000000000000000007465207263746F20313230",
      INIT_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_07 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_08 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_09 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_0F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 256 to 511, Port B Address 128 to 255
      INIT_10 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_11 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_12 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_13 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_14 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_15 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_16 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_17 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_18 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_19 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_1F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 512 to 767, Port B Address 256 to 383
      INIT_20 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_21 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_22 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_23 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_24 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_25 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_26 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_27 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_28 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_29 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_2F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 768 to 1023, Port B Address 384 to 511
      INIT_30 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_31 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_32 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_33 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_34 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_35 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_36 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_37 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_38 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_39 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3A => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3B => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3C => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3D => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3E => X"0000000000000000000000000000000000000000000000000000000000000000",
      INIT_3F => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- The next set of INITP_xx are for the parity bits
      -- Port A Address 0 to 255, Port B Address 0 to 127
      INITP_00 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_01 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 256 to 511, Port B Address 128 to 255
      INITP_02 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_03 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 512 to 767, Port B Address 256 to 383
      INITP_04 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_05 => X"0000000000000000000000000000000000000000000000000000000000000000",
      -- Port A Address 768 to 1023, Port B Address 384 to 511
      INITP_06 => X"0000000000000000000000000000000000000000000000000000000000000000",
      INITP_07 => X"0000000000000000000000000000000000000000000000000000000000000000")
   port map (
      DOA => open,--DOA,    --  DOA,      -- Port A 16-bit Data Output
      DOB => D(16-1 downto 8),--D(8-1 downto 0),--DOB,      -- Port B 8-bit Data Output
      DOPA => open,--DOPA,    -- Port A 2-bit Parity Output
      DOPB => open,--DOPB,    -- Port B 1-bit Parity Output
      ADDRA => "0000000000",--A,  --  ADDRA,  -- Port A 10-bit Address Input
      ADDRB => ADDRB,  -- Port B 11-bit Address Input
      CLKA => '0',--Clk, --  CLKA,    -- Port A 1-bit Clock
      CLKB => Clk,--CLKB,    -- Port B 1-bit Clock
      DIA => DIA,      -- Port A 16-bit Data Input
      DIB => DIB,      -- Port B 8-bit Data Input
      DIPA => DIPA,    -- Port A 2-bit parity Input
      DIPB => DIPB,    -- Port B 1-bit parity Input
      ENA => ENA,      -- Port A 1-bit RAM Enable Input
      ENB => '1',--ENB,      -- Port B 1-bit RAM Enable Input
      SSRA => SSRA,    -- Port A 1-bit Synchronous Set/Reset Input
      SSRB => SSRB,    -- Port B 1-bit Synchronous Set/Reset Input
      WEA => WEA,      -- Port A 2-bit Write Enable Input
      WEB => WEB       -- Port B 1-bit Write Enable Input
   );

end Behavioral;

