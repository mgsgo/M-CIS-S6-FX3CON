# This file was generated with hex2rom written by Daniel Wallner

INST *brom231300 INIT_00 = 1D01B0A610D1B1A60D31C803F1ECB0A010CDCF1F111A1B1C221E1F202122230A;
INST *brom231300 INIT_01 = 8CFE5F08899A98181F0F0F0F8F86808C8F110F0F0F1F088CFE5DDA8768E1B1A8;
INST *brom231300 INIT_02 = 08EFFF0F1FCFDFACDFCE21D1901F0E81F1E008D0C01908F7E6DFCF1F0FFFEF08;
INST *brom231300 INIT_03 = 09F1E0908D298A80FFEE2109F1E0900F1006DFCEF9FDECDFCEE8DFCF1F0FFFEF;
INST *brom231300 INIT_04 = 88868078C49087A870669080898A8A8882818FF808EFFF0F1FCFDF618888FDEC;
INST *brom231300 INIT_05 = 74697465207263746F20313230540020534DFFF8F19695A180F6961189FA9511;
INST *brom231300 INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000;
INST *brom231301 INIT_00 = 92C0E0E8E0F70738929695C0E0E5E0E6E0BFEDBE24C0C0C0C0C0C0C0C0C0C0C0;
INST *brom231301 INIT_01 = B1CF9B95B9B9E9959090BE90910093B1932492B6929295B9CF9BCFC0D0F70738;
INST *brom231301 INIT_02 = 95909091919191F3051596DFE02F2F912F2FC0E0E02F2F2E2E93939393929295;
INST *brom231301 INIT_03 = 952F2FE0E0F430812D2D96952F2FE0C0E0E22D2D2E2E2E2D2D2E939393939292;
INST *brom231301 INIT_04 = 33009194DFE0E6DFE0E0E0E6B9E1B9E9BBBBEF9495909091919191F723812E2E;
INST *brom231301 INIT_05 = 006E207374656F20667333335339410A4747CF94CF9898F733CF9AF433CF9AF4;
INST *brom231301 INIT_06 = 0000000000000000000000000000000000000000000000000000000000000000;
